`include "A4Q1_fsm.v"

module tb();
    reg in;
    reg [2:0] state;
    wire out;

    fsm
endmodule