module fsm_driver()