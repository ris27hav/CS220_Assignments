`include "A4Q1_fsm_driver.v"

module tb();
    reg in;
    reg [2:0] state;
    wire out;

    fsm
endmodule