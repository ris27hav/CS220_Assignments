`include "A4Q1_fsm.v"

module tb();
    reg [7:0] in;
    reg [2:0] state;
    wire [7:0] out;

    fsm
endmodule